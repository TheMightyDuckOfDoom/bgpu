// Copyright 2025 Tobias Senti
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51

`ifndef BGPU_INSTRUCTIONS_SVH_
`define BGPU_INSTRUCTIONS_SVH_

typedef enum logic [1:0] {
    BGPU_EU_IU  = 'd0,
    BGPU_EU_LSU = 'd1
} bgpu_eu_e;

typedef enum logic [5:0] {
    IU_TID  = 'h00, // Get thread ID inside a warp
    IU_WID  = 'h01, // Get warp ID

    IU_ADD  = 'h02, // Add operands
    IU_SUB  = 'h03, // Subtract operands
    IU_AND  = 'h04, // Bitwise AND operands
    IU_OR   = 'h05, // Bitwise OR operands
    IU_XOR  = 'h06, // Bitwise XOR operands

    IU_LDI  = 'h07, // Load immediate -> concatenate operands register index
    IU_ADDI = 'h08, // Add immediate -> add immediate value to first operand
    IU_SUBI = 'h09, // Subtract immediate -> subtract immediate value from first operand

    IU_SLL  = 'h0A, // Shift left logical
    IU_SLLI = 'h0B  // Shift left logical immediate
} bgpu_iu_subtype_e;

typedef enum logic [5:0] {
    LSU_LOAD_BYTE  = 'h00, // Load from memory
    LSU_LOAD_HALF  = 'h01, // Load half-word from memory
    LSU_LOAD_WORD  = 'h02, // Load word from memory
    LSU_STORE_BYTE = 'h03, // Store byte to memory
    LSU_STORE_HALF = 'h04, // Store half-word to memory
    LSU_STORE_WORD = 'h05  // Store word to memory
} bgpu_lsu_subtype_e;

typedef union packed {
    bgpu_iu_subtype_e  iu;
    bgpu_lsu_subtype_e lsu;
} bgpu_inst_subtype_u;

typedef struct packed {
    bgpu_eu_e           eu;
    bgpu_inst_subtype_u subtype;
} bgpu_inst_t;

// Both operands are registers
`define BGPU_IU_TWO_REG_OPERANDS {\
    IU_ADD,\
    IU_SUB,\
    IU_AND,\
    IU_OR,\
    IU_XOR,\
    IU_SLL\
}

// First operand is an immediate, second is an register
`define BGPU_IU_REG_IMM_OPERANDS {\
    IU_ADDI,\
    IU_SUBI,\
    IU_SLLI\
}

// Store operations
`define BGPU_INST_STORE {\
    LSU_STORE_BYTE,\
    LSU_STORE_HALF,\
    LSU_STORE_WORD\
}

`define BGPU_INST_LOAD {\
    LSU_LOAD_BYTE,\
    LSU_LOAD_HALF,\
    LSU_LOAD_WORD\
}

`ifndef SYNTHESIS
    `define BGPU_INT_UNIT_VALID_SUBTYPES {\
        IU_TID,\
        IU_WID,\
        IU_ADD,\
        IU_SUB,\
        IU_AND,\
        IU_OR,\
        IU_XOR,\
        IU_LDI,\
        IU_ADDI,\
        IU_SUBI,\
        IU_SLL,\
        IU_SLLI\
    }
`endif

`endif
