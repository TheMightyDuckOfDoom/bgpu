// Copyright 2025 Tobias Senti
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51

/// Compute Unit
module compute_unit import bgpu_pkg::*; #(
    /// Width of the Program Counter
    parameter int unsigned PcWidth = 16,
    /// Number of warps
    parameter int unsigned NumWarps = 8,
    /// Number of threads per warp
    parameter int unsigned WarpWidth = 4,
    /// Encoded instruction width
    parameter int unsigned EncInstWidth = 32,
    /// Number of inflight instructions per warp
    parameter int unsigned InflightInstrPerWarp = 4,
    /// How many registers can each warp access as operand or destination
    parameter int unsigned RegIdxWidth = 8,
    /// How many operands each instruction can have
    parameter int unsigned OperandsPerInst = 2,
    /// How many register banks are available
    parameter int unsigned NumBanks = 4,
    /// How many operand collectors are available
    parameter int unsigned NumOperandCollectors = 6,
    /// Should the register banks be dual ported?
    parameter bit          DualPortRegisterBanks = 1'b0,
    /// Width of the registers
    parameter int unsigned RegWidth = 32,
    // Memory Address width in bits
    parameter int unsigned AddressWidth = 32,
    // Memory Block size in bytes -> Memory request width
    parameter int unsigned BlockIdxBits = 4,
    // Width of the id for requests queue
    parameter int unsigned OutstandingReqIdxWidth = 3,
    // Number of cache lines in the instruction cache
    parameter int unsigned NumIClines = 8,
    // Number of bits for the instruction cache line index
    parameter int unsigned IClineIdxBits = 2,
    // How many bits are used to index thread blocks inside a thread group?
    parameter int unsigned TblockIdxBits = 8,
    // How many bits are used to identify a thread block?
    parameter int unsigned TblockIdBits = 8,

    /// Dependent parameter, do **not** overwrite.
    parameter int unsigned BlockAddrWidth  = AddressWidth - BlockIdxBits,
    parameter int unsigned BlockWidth      = 1 << BlockIdxBits, // In bytes
    parameter int unsigned ThreadIdxWidth  = WarpWidth > 1 ? $clog2(WarpWidth) : 1,
    parameter int unsigned ICAddrWidth     = IClineIdxBits > 0 ? PcWidth - IClineIdxBits : PcWidth,
    parameter type tblock_idx_t = logic      [       TblockIdxBits-1:0],
    parameter type tblock_id_t  = logic      [        TblockIdBits-1:0],
    parameter type addr_t       = logic      [        AddressWidth-1:0],
    parameter type imem_addr_t  = logic      [         ICAddrWidth-1:0],
    parameter type enc_inst_t   = logic      [        EncInstWidth-1:0],
    parameter type imem_data_t  = enc_inst_t [(1 << IClineIdxBits)-1:0],
    parameter type pc_t         = logic      [             PcWidth-1:0],
    parameter type block_addr_t = logic      [      BlockAddrWidth-1:0],
    parameter type byte_t       = logic      [                     7:0],
    parameter type block_data_t = byte_t     [          BlockWidth-1:0],
    parameter type block_idx_t  = logic      [        BlockIdxBits-1:0],
    parameter type block_mask_t = logic      [          BlockWidth-1:0],
    parameter type req_id_t     = logic      [OutstandingReqIdxWidth + ThreadIdxWidth-1:0]
) (
    // Clock and reset
    input logic clk_i,
    input logic rst_ni,

    // Interface to start a new thread block on this compute unit
    output logic        warp_free_o, // The is atleas one free warp that can start a new block
    input  logic        allocate_warp_i,
    input  pc_t         allocate_pc_i,
    input  addr_t       allocate_dp_addr_i, // Data / Parameter address
    input  tblock_idx_t allocate_tblock_idx_i, // Block index -> used to calculate the thread id
    input  tblock_id_t  allocate_tblock_id_i,  // Block id -> unique identifier for the block

    // Thread block completion
    output logic       tblock_done_o,
    output tblock_id_t tblock_done_id_o,

    /// Instruction Memory Request
    input  logic       imem_ready_i,
    output logic       imem_req_valid_o,
    output imem_addr_t imem_req_addr_o,

    /// Instruction Memory Response
    input  logic       imem_rsp_valid_i,
    input  imem_data_t imem_rsp_data_i,

    /// Memory Request
    input  logic        mem_ready_i,
    output logic        mem_req_valid_o,
    output req_id_t     mem_req_id_o,
    output block_addr_t mem_req_addr_o,
    output block_mask_t mem_req_we_mask_o,
    output block_data_t mem_req_wdata_o,

    /// Memory Response
    input  logic        mem_rsp_valid_i,
    input  req_id_t     mem_rsp_id_i,
    input  block_data_t mem_rsp_data_i
);
    // #######################################################################################
    // # Local Parameters                                                                    #
    // #######################################################################################

    localparam int unsigned NumTags  = InflightInstrPerWarp;
    localparam int unsigned WidWidth = NumWarps > 1 ? $clog2(NumWarps) : 1;
    localparam int unsigned TagWidth = NumTags > 1  ? $clog2(NumTags)  : 1;

    // #######################################################################################
    // # Typedefs                                                                            #
    // #######################################################################################

    // Typedefs
    typedef logic [         RegIdxWidth-1:0] reg_idx_t;
    typedef logic [ WidWidth + TagWidth-1:0] iid_t;
    typedef logic [           WarpWidth-1:0] act_mask_t;
    typedef logic [RegWidth * WarpWidth-1:0] warp_data_t;
    typedef logic [    WidWidth-1:0] wid_t;

    // Fetcher to Instruction Cache type
    typedef struct packed {
        pc_t       pc;
        act_mask_t act_mask;
        wid_t      warp_id;
    } fe_to_ic_data_t;

    // Instruction Cache to Decoder type
    typedef struct packed {
        pc_t       pc;
        act_mask_t act_mask;
        wid_t      warp_id;
        enc_inst_t inst;
    } ic_to_dec_data_t;

    // Decoder to Instruction Buffer type
    typedef struct packed {
        pc_t       pc;
        act_mask_t act_mask;
        wid_t      warp_id;
        inst_t     inst;
        reg_idx_t  dst;
        logic      [OperandsPerInst-1:0] operands_required;
        reg_idx_t  [OperandsPerInst-1:0] operands;
    } dec_to_ib_data_t;

    // Multi Warp Dispatcher to Register Operand Collector Stage type
    typedef struct packed {
        iid_t      tag;
        pc_t       pc;
        act_mask_t act_mask;
        inst_t     inst;
        reg_idx_t  dst;
        logic      [OperandsPerInst-1:0] operands_required;
        reg_idx_t  [OperandsPerInst-1:0] operands;
    } disp_to_opc_data_t;

    // Register Operand Collector Stage to Execution Units type
    typedef struct packed {
        iid_t       tag;
        pc_t        pc;
        act_mask_t  act_mask;
        inst_t      inst;
        reg_idx_t   dst;
        warp_data_t [OperandsPerInst-1:0] operands;
    } opc_to_eu_data_t;

    // Execution Units to Register Operand Collector Stage type
    typedef struct packed {
        iid_t       tag;
        reg_idx_t   dst;
        warp_data_t data;
    } eu_to_opc_data_t;

    // #######################################################################################
    // # Signals                                                                             #
    // #######################################################################################


    // Fetcher to Instruction Cache
    logic fe_to_ic_valid_d, fe_to_ic_valid_q;
    logic ic_to_fe_ready_d, ic_to_fe_ready_q;
    fe_to_ic_data_t fe_to_ic_data_d, fe_to_ic_data_q;

    // Fetcher to Integer Unit -> Constants per Warp
    addr_t       [NumWarps-1:0] fe_to_iu_warp_dp_addr;    // Data / Parameter address
    tblock_idx_t [NumWarps-1:0] fe_to_iu_warp_tblock_idx; // Block index

    /// Instruction Cache to Decoder
    logic ic_to_dec_valid, dec_to_ic_ready;
    ic_to_dec_data_t ic_to_dec_data;

    // Decoder to Fetcher
    logic dec_to_fetch_decoded;
    logic dec_to_fetch_stop_warp;
    wid_t dec_to_fetch_decoded_warp_id;
    pc_t  dec_to_fetch_decoded_next_pc;

    // Decoder to Instruction Buffer
    logic dec_to_ib_valid_d, dec_to_ib_valid_q;
    logic ib_to_dec_ready_d, ib_to_dec_ready_q;
    dec_to_ib_data_t dec_to_ib_data_d, dec_to_ib_data_q;

    // Instruction Buffer to Fetcher
    logic [NumWarps-1:0] ib_space_available; // Which warp has space for a new instruction?
    logic [NumWarps-1:0] ib_all_instr_finished; // Are there any instructions in flight?

    // Multi Warp Dispatcher to Register Operand Collector Stage
    logic disp_to_opc_valid, opc_to_disp_ready;
    disp_to_opc_data_t disp_to_opc_data;

    // Register Operand Collector Stage to Execution Units
    logic opc_to_eu_valid,  eu_to_opc_ready;
    logic opc_to_iu_valid,  iu_to_opc_ready;
    logic opc_to_lsu_valid, lsu_to_opc_ready;
    opc_to_eu_data_t opc_to_eu_data;

    // Execution Units to Register Operand Collector Stage
    logic eu_to_opc_valid, opc_to_eu_ready;
    logic iu_to_rc_valid,  rc_to_iu_ready;
    logic lsu_to_rc_valid, rc_to_lsu_ready;
    eu_to_opc_data_t eu_to_opc_data, iu_to_rc_data, lsu_to_rc_data;

    // #######################################################################################
    // # Fetcher                                                                             #
    // #######################################################################################

    fetcher #(
        .PcWidth      ( PcWidth       ),
        .NumWarps     ( NumWarps      ),
        .WarpWidth    ( WarpWidth     ),
        .AddressWidth ( AddressWidth  ),
        .TblockIdxBits( TblockIdxBits ),
        .TblockIdBits ( TblockIdBits  )
    ) i_fetcher (
        .clk_i ( clk_i  ),
        .rst_ni( rst_ni ),

        .warp_free_o          ( warp_free_o           ),
        .allocate_warp_i      ( allocate_warp_i       ),
        .allocate_pc_i        ( allocate_pc_i         ),
        .allocate_dp_addr_i   ( allocate_dp_addr_i    ),
        .allocate_tblock_idx_i( allocate_tblock_idx_i ),
        .allocate_tblock_id_i ( allocate_tblock_id_i  ),

        .tblock_done_o   ( tblock_done_o    ),
        .tblock_done_id_o( tblock_done_id_o ),

        .ib_space_available_i   ( ib_space_available    ),
        .ib_all_instr_finished_i( ib_all_instr_finished ),

        .ic_ready_i   ( ic_to_fe_ready_q         ),
        .fe_valid_o   ( fe_to_ic_valid_d         ),
        .fe_pc_o      ( fe_to_ic_data_d.pc       ),
        .fe_act_mask_o( fe_to_ic_data_d.act_mask ),
        .fe_warp_id_o ( fe_to_ic_data_d.warp_id  ),

        .dec_decoded_i        ( dec_to_fetch_decoded         ),
        .dec_stop_warp_i      ( dec_to_fetch_stop_warp       ),
        .dec_decoded_warp_id_i( dec_to_fetch_decoded_warp_id ),
        .dec_decoded_next_pc_i( dec_to_fetch_decoded_next_pc ),

        .warp_dp_addr_o   ( fe_to_iu_warp_dp_addr    ),
        .warp_tblock_idx_o( fe_to_iu_warp_tblock_idx )
    );

    // #######################################################################################
    // # Fetcher to Instruction Cache - Register                                             #
    // #######################################################################################

    stream_register #(
        .T( fe_to_ic_data_t )
    ) i_fe_to_ic_reg (
        .clk_i     ( clk_i  ),
        .rst_ni    ( rst_ni ),
        .clr_i     ( 1'b0   ),
        .testmode_i( 1'b0   ),

        .valid_i( fe_to_ic_valid_d ),
        .ready_o( ic_to_fe_ready_q ),
        .data_i ( fe_to_ic_data_d  ),

        .valid_o( fe_to_ic_valid_q ),
        .ready_i( ic_to_fe_ready_d ),
        .data_o ( fe_to_ic_data_q  )
    );

    // #######################################################################################
    // # Instruction Cache                                                                   #
    // #######################################################################################

    instruction_cache #(
        .PcWidth         ( PcWidth       ),
        .NumWarps        ( NumWarps      ),
        .WarpWidth       ( WarpWidth     ),
        .EncInstWidth    ( EncInstWidth  ),
        .CachelineIdxBits( IClineIdxBits ),
        .NumCachelines   ( NumIClines    )
    ) i_instruction_cache (
        .clk_i ( clk_i  ),
        .rst_ni( rst_ni ),

        .mem_ready_i( imem_ready_i     ),
        .mem_req_o  ( imem_req_valid_o ),
        .mem_addr_o ( imem_req_addr_o  ),

        .mem_valid_i( imem_rsp_valid_i ),
        .mem_data_i ( imem_rsp_data_i  ),

        .ic_ready_o   ( ic_to_fe_ready_d         ),
        .fe_valid_i   ( fe_to_ic_valid_q         ),
        .fe_pc_i      ( fe_to_ic_data_q.pc       ),
        .fe_act_mask_i( fe_to_ic_data_q.act_mask ),
        .fe_warp_id_i ( fe_to_ic_data_q.warp_id  ),

        .dec_ready_i  ( dec_to_ic_ready         ),
        .ic_valid_o   ( ic_to_dec_valid         ),
        .ic_pc_o      ( ic_to_dec_data.pc       ),
        .ic_act_mask_o( ic_to_dec_data.act_mask ),
        .ic_warp_id_o ( ic_to_dec_data.warp_id  ),
        .ic_inst_o    ( ic_to_dec_data.inst     )
    );

    // #######################################################################################
    // # Instruction Decoder                                                                 #
    // #######################################################################################

    decoder #(
        .PcWidth        ( PcWidth         ),
        .NumWarps       ( NumWarps        ),
        .WarpWidth      ( WarpWidth       ),
        .EncInstWidth   ( EncInstWidth    ),
        .RegIdxWidth    ( RegIdxWidth     ),
        .OperandsPerInst( OperandsPerInst )
    ) i_decoder (
        .dec_ready_o  ( dec_to_ic_ready         ),
        .ic_valid_i   ( ic_to_dec_valid         ),
        .ic_pc_i      ( ic_to_dec_data.pc       ),
        .ic_act_mask_i( ic_to_dec_data.act_mask ),
        .ic_warp_id_i ( ic_to_dec_data.warp_id  ),
        .ic_inst_i    ( ic_to_dec_data.inst     ),

        .disp_ready_i           ( ib_to_dec_ready_q                  ),
        .dec_valid_o            ( dec_to_ib_valid_d                  ),
        .dec_pc_o               ( dec_to_ib_data_d.pc                ),
        .dec_act_mask_o         ( dec_to_ib_data_d.act_mask          ),
        .dec_warp_id_o          ( dec_to_ib_data_d.warp_id           ),
        .dec_inst_o             ( dec_to_ib_data_d.inst              ),
        .dec_dst_o              ( dec_to_ib_data_d.dst               ),
        .dec_operands_required_o( dec_to_ib_data_d.operands_required ),
        .dec_operands_o         ( dec_to_ib_data_d.operands          ),

        .dec_decoded_o         ( dec_to_fetch_decoded         ),
        .dec_stop_warp_o       ( dec_to_fetch_stop_warp       ),
        .dec_decoded_warp_id_o ( dec_to_fetch_decoded_warp_id ),
        .dec_decoded_next_pc_o ( dec_to_fetch_decoded_next_pc )
    );

    // #######################################################################################
    // # Decoder to Instruction Buffer - Register                                            #
    // #######################################################################################

    stream_register #(
        .T( dec_to_ib_data_t )
    ) i_dec_to_ib_reg (
        .clk_i     ( clk_i  ),
        .rst_ni    ( rst_ni ),
        .clr_i     ( 1'b0   ),
        .testmode_i( 1'b0   ),

        .valid_i( dec_to_ib_valid_d ),
        .ready_o( ib_to_dec_ready_q ),
        .data_i ( dec_to_ib_data_d  ),

        .valid_o( dec_to_ib_valid_q ),
        .ready_i( ib_to_dec_ready_d ),
        .data_o ( dec_to_ib_data_q  )
    );

    // #######################################################################################
    // # Multi Warp Dispatcher                                                               #
    // #######################################################################################

    multi_warp_dispatcher #(
        .NumTags              ( NumTags               ),
        .PcWidth              ( PcWidth               ),
        .NumWarps             ( NumWarps              ),
        .WarpWidth            ( WarpWidth             ),
        .WaitBufferSizePerWarp( InflightInstrPerWarp  ),
        .RegIdxWidth          ( RegIdxWidth           ),
        .OperandsPerInst      ( OperandsPerInst       )
    ) i_warp_dispatcher (
        .clk_i ( clk_i  ),
        .rst_ni( rst_ni ),

        .fe_handshake_i( fe_to_ic_valid_d && ic_to_fe_ready_q ),
        .fe_warp_id_i  ( fe_to_ic_data_d.warp_id              ),

        .ib_space_available_o   ( ib_space_available    ),
        .ib_all_instr_finished_o( ib_all_instr_finished ),

        .dec_stop_decoded_i        ( dec_to_fetch_decoded && dec_to_fetch_stop_warp ),
        .dec_stop_decoded_warp_id_i( dec_to_fetch_decoded_warp_id                   ),

        .ib_ready_o             ( ib_to_dec_ready_d                  ),
        .dec_valid_i            ( dec_to_ib_valid_q                  ),
        .dec_pc_i               ( dec_to_ib_data_q.pc                ),
        .dec_act_mask_i         ( dec_to_ib_data_q.act_mask          ),
        .dec_warp_id_i          ( dec_to_ib_data_q.warp_id           ),
        .dec_inst_i             ( dec_to_ib_data_q.inst              ),
        .dec_dst_i              ( dec_to_ib_data_q.dst               ),
        .dec_operands_required_i( dec_to_ib_data_q.operands_required ),
        .dec_operands_i         ( dec_to_ib_data_q.operands          ),

        .opc_ready_i             ( opc_to_disp_ready                  ),
        .disp_valid_o            ( disp_to_opc_valid                  ),
        .disp_tag_o              ( disp_to_opc_data.tag               ),
        .disp_pc_o               ( disp_to_opc_data.pc                ),
        .disp_act_mask_o         ( disp_to_opc_data.act_mask          ),
        .disp_inst_o             ( disp_to_opc_data.inst              ),
        .disp_dst_o              ( disp_to_opc_data.dst               ),
        .disp_operands_required_o( disp_to_opc_data.operands_required ),
        .disp_operands_o         ( disp_to_opc_data.operands          ),

        .eu_valid_i( eu_to_opc_valid && opc_to_eu_ready ),
        .eu_tag_i  ( eu_to_opc_data.tag                 )
    );

    // #######################################################################################
    // # Register Operand Collector Stage                                                    #
    // #######################################################################################

    register_opc_stage #(
        .NumTags              ( NumTags               ),
        .PcWidth              ( PcWidth               ),
        .NumWarps             ( NumWarps              ),
        .WarpWidth            ( WarpWidth             ),
        .RegIdxWidth          ( RegIdxWidth           ),
        .OperandsPerInst      ( OperandsPerInst       ),
        .NumBanks             ( NumBanks              ),
        .RegWidth             ( RegWidth              ),
        .DualPortRegisterBanks( DualPortRegisterBanks ),
        .NumOperandCollectors ( NumOperandCollectors  )
    ) i_register_opc_stage (
        .clk_i ( clk_i  ),
        .rst_ni( rst_ni ),

        .opc_ready_o        ( opc_to_disp_ready                  ),
        .disp_valid_i       ( disp_to_opc_valid                  ),
        .disp_tag_i         ( disp_to_opc_data.tag               ),
        .disp_pc_i          ( disp_to_opc_data.pc                ),
        .disp_act_mask_i    ( disp_to_opc_data.act_mask          ),
        .disp_inst_i        ( disp_to_opc_data.inst              ),
        .disp_dst_i         ( disp_to_opc_data.dst               ),
        .disp_src_required_i( disp_to_opc_data.operands_required ),
        .disp_src_i         ( disp_to_opc_data.operands          ),

        .eu_ready_i        ( eu_to_opc_ready         ),
        .opc_valid_o       ( opc_to_eu_valid         ),
        .opc_tag_o         ( opc_to_eu_data.tag      ),
        .opc_pc_o          ( opc_to_eu_data.pc       ),
        .opc_act_mask_o    ( opc_to_eu_data.act_mask ),
        .opc_inst_o        ( opc_to_eu_data.inst     ),
        .opc_dst_o         ( opc_to_eu_data.dst      ),
        .opc_operand_data_o( opc_to_eu_data.operands ),

        .opc_to_eu_ready_o( opc_to_eu_ready     ),
        .eu_valid_i       ( eu_to_opc_valid     ),
        .eu_tag_i         ( eu_to_opc_data.tag  ),
        .eu_dst_i         ( eu_to_opc_data.dst  ),
        .eu_data_i        ( eu_to_opc_data.data )
    );

    // #######################################################################################
    // # Execution Unit Demux                                                                #
    // #######################################################################################

    stream_demux #(
        .N_OUP(2)
    ) i_eu_demux (
        .inp_valid_i( opc_to_eu_valid ),
        .inp_ready_o( eu_to_opc_ready ),

        .oup_sel_i( opc_to_eu_data.inst.eu[0] ),

        .oup_valid_o({ opc_to_lsu_valid, opc_to_iu_valid }),
        .oup_ready_i({ lsu_to_opc_ready, iu_to_opc_ready })
    );

    `ifndef SYNTHESIS
        assert property (@(posedge clk_i) opc_to_eu_valid
            |-> opc_to_eu_data.inst.eu inside {EU_IU, EU_LSU})
            else $error("Invalid execution unit type: %0d", opc_to_eu_data.inst.eu);
    `endif

    // #######################################################################################
    // # Execution Units                                                                     #
    // #######################################################################################

    // Integer Unit
    integer_unit #(
        .NumTags        ( NumTags         ),
        .NumWarps       ( NumWarps        ),
        .RegWidth       ( RegWidth        ),
        .WarpWidth      ( WarpWidth       ),
        .OperandsPerInst( OperandsPerInst ),
        .RegIdxWidth    ( RegIdxWidth     ),
        .AddressWidth   ( AddressWidth    ),
        .TblockIdxBits  ( TblockIdxBits   )
    ) i_integer_unit (
        .clk_i ( clk_i  ),
        .rst_ni( rst_ni ),

        .fe_to_iu_warp_dp_addr_i   ( fe_to_iu_warp_dp_addr    ),
        .fe_to_iu_warp_tblock_idx_i( fe_to_iu_warp_tblock_idx ),

        .eu_to_opc_ready_o   ( iu_to_opc_ready                ),
        .opc_to_eu_valid_i   ( opc_to_iu_valid                ),
        .opc_to_eu_tag_i     ( opc_to_eu_data.tag             ),
        .opc_to_eu_inst_sub_i( opc_to_eu_data.inst.subtype.iu ),
        .opc_to_eu_dst_i     ( opc_to_eu_data.dst             ),
        .opc_to_eu_operands_i( opc_to_eu_data.operands        ),

        .rc_to_eu_ready_i( rc_to_iu_ready     ),
        .eu_to_rc_valid_o( iu_to_rc_valid     ),
        .eu_to_rc_tag_o  ( iu_to_rc_data.tag  ),
        .eu_to_rc_dst_o  ( iu_to_rc_data.dst  ),
        .eu_to_rc_data_o ( iu_to_rc_data.data )
    );

    // Load Store Unit
    load_store_unit #(
        .RegWidth              ( RegWidth               ),
        .WarpWidth             ( WarpWidth              ),
        .OperandsPerInst       ( OperandsPerInst        ),
        .RegIdxWidth           ( RegIdxWidth            ),
        .iid_t                 ( iid_t                  ),
        .AddressWidth          ( AddressWidth           ),
        .BlockIdxBits          ( BlockIdxBits           ),
        .OutstandingReqIdxWidth( OutstandingReqIdxWidth )
    ) i_load_store_unit (
        .clk_i ( clk_i  ),
        .rst_ni( rst_ni ),

        .eu_to_opc_ready_o   ( lsu_to_opc_ready                ),
        .opc_to_eu_valid_i   ( opc_to_lsu_valid                ),
        .opc_to_eu_tag_i     ( opc_to_eu_data.tag              ),
        .opc_to_eu_inst_sub_i( opc_to_eu_data.inst.subtype.lsu ),
        .opc_to_eu_act_mask_i( opc_to_eu_data.act_mask         ),
        .opc_to_eu_dst_i     ( opc_to_eu_data.dst              ),
        .opc_to_eu_operands_i( opc_to_eu_data.operands         ),

        .rc_to_eu_ready_i( rc_to_lsu_ready     ),
        .eu_to_rc_valid_o( lsu_to_rc_valid     ),
        .eu_to_rc_tag_o  ( lsu_to_rc_data.tag  ),
        .eu_to_rc_dst_o  ( lsu_to_rc_data.dst  ),
        .eu_to_rc_data_o ( lsu_to_rc_data.data ),

        .mem_ready_i      ( mem_ready_i       ),
        .mem_req_valid_o  ( mem_req_valid_o   ),
        .mem_req_id_o     ( mem_req_id_o      ),
        .mem_req_addr_o   ( mem_req_addr_o    ),
        .mem_req_we_mask_o( mem_req_we_mask_o ),
        .mem_req_wdata_o  ( mem_req_wdata_o   ),

        .mem_rsp_valid_i  ( mem_rsp_valid_i   ),
        .mem_rsp_id_i     ( mem_rsp_id_i      ),
        .mem_rsp_data_i   ( mem_rsp_data_i    )
    );

    // #######################################################################################
    // # Execution Unit Result Collector                                                     #
    // #######################################################################################

    stream_arbiter #(
        .DATA_T ( eu_to_opc_data_t ),
        .N_INP  ( 2                ),
        .ARBITER( "rr"             )
    ) i_result_collector (
        .clk_i        ( clk_i           ),
        .rst_ni       ( rst_ni          ),
        .inp_data_i   ({ iu_to_rc_data,  lsu_to_rc_data  }),
        .inp_valid_i  ({ iu_to_rc_valid, lsu_to_rc_valid }),
        .inp_ready_o  ({ rc_to_iu_ready, rc_to_lsu_ready }),

        .oup_data_o   ( eu_to_opc_data   ),
        .oup_valid_o  ( eu_to_opc_valid  ),
        .oup_ready_i  ( opc_to_eu_ready  )
    );

endmodule : compute_unit
